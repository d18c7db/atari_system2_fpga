--	(c) 2020 d18c7db(a)hotmail
--
--	This program is free software; you can redistribute it and/or modify it under
--	the terms of the GNU General Public License version 3 or, at your option,
--	any later version as published by the Free Software Foundation.
--
--	This program is distributed in the hope that it will be useful,
--	but WITHOUT ANY WARRANTY; without even the implied warranty of
--	MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.
--
-- For full details, see the GNU General Public License at www.gnu.org/licenses
--
-- generic 2K x 8 RAM definition

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;

entity RAM_8K16 is
	port(
		I_MCKR : in  std_logic;
		I_En   : in  std_logic;
		I_Wn   : in  std_logic;
		I_ADDR : in  std_logic_vector(12 downto 0);
		I_DATA : in  std_logic_vector(15 downto 0);
		O_DATA : out std_logic_vector(15 downto 0)
	);
end RAM_8K16;

architecture RTL of RAM_8K16 is
	type RAM_ARRAY_8Kx16 is array (0 to 8191) of std_logic_vector(15 downto 0);
	signal RAM : RAM_ARRAY_8Kx16 := (
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F00", x"1F00", x"1F00", x"1F00", x"1F00", x"1F00",
	x"1F00", x"1F00", x"1F00", x"1F00", x"1F00", x"1F00", x"1F00", x"1F00",
	x"1F00", x"1F00", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F00", x"1F00", x"1F00", x"1F00", x"1F00", x"1F02",
	x"1F03", x"1F04", x"1F00", x"1F00", x"1F00", x"1F00", x"1F05", x"1F06",
	x"1F11", x"1F12", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F00", x"1F00", x"1F00", x"1F18", x"1F13", x"1F14",
	x"1F15", x"1F16", x"1F17", x"1F1C", x"1F00", x"1F1D", x"1F1E", x"1F1F",
	x"1F20", x"1F21", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F00", x"1F00", x"1F00", x"1F22", x"1F23", x"1F24",
	x"1F25", x"1F26", x"1F27", x"1F28", x"1F2B", x"1F2C", x"1F2D", x"1F2E",
	x"1F2F", x"1F30", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F00", x"1F00", x"1F31", x"1F32", x"1F33", x"1F34",
	x"1F35", x"1F36", x"1F37", x"1F38", x"1F39", x"1F3A", x"1F3B", x"1F3C",
	x"1F3D", x"1F3E", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F00", x"1F00", x"1F3F", x"1F40", x"1F41", x"1F42",
	x"1F43", x"1F44", x"1F45", x"1F46", x"1F47", x"1F48", x"1F49", x"1F4A",
	x"1F4B", x"1F4C", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F00", x"1F00", x"1F4D", x"1F4E", x"1F4F", x"1F50",
	x"1F51", x"1F52", x"1F53", x"1F54", x"1F55", x"1F56", x"1F57", x"1F58",
	x"1F59", x"1F5A", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F00", x"1F5B", x"1F5C", x"1F5D", x"1F5E", x"1F5F",
	x"1F60", x"1F61", x"1F62", x"1F63", x"1F64", x"1F65", x"1F66", x"1F67",
	x"1F68", x"1F00", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F69", x"1F6A", x"1F6B", x"1F6C", x"1F6D", x"1F6E",
	x"1F6F", x"1F70", x"1F71", x"1F72", x"1F73", x"1F74", x"1F75", x"1F76",
	x"1F77", x"1F00", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F78", x"1F79", x"1F7A", x"1F7B", x"1F7C", x"1F7D",
	x"1F7E", x"1F81", x"1F82", x"1F83", x"1F84", x"1F85", x"1F86", x"1F87",
	x"1F88", x"1F89", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F8A", x"1F8B", x"1F8C", x"1F8D", x"1F8E", x"1F8F",
	x"1F90", x"1F91", x"1F92", x"1F93", x"1F00", x"1F94", x"1F95", x"1F96",
	x"1F97", x"1F98", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F99", x"1F00", x"1F00", x"1F9A", x"1F9B", x"1F9C",
	x"1F9D", x"1F9E", x"1F9F", x"1FA0", x"1FA1", x"1FA2", x"1FA3", x"1FA4",
	x"1FA5", x"1FA6", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F00", x"1F00", x"1FA7", x"1FA8", x"1FA9", x"1FAA",
	x"1FAB", x"1FAC", x"1FAD", x"1FAE", x"1FAF", x"1FB0", x"1FB1", x"1FB2",
	x"1FB3", x"1FB4", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1F00", x"1FB5", x"1FB6", x"1FB7", x"1FB8", x"1FB9",
	x"1FBA", x"1FBB", x"1FBC", x"1FBD", x"1FBE", x"1FBF", x"1FC0", x"1FC1",
	x"1FC2", x"1FC3", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1FC4", x"1FC5", x"1FC6", x"1FC7", x"1FC8", x"1FC9",
	x"1FCA", x"1FCB", x"1FCC", x"1FCD", x"1FCE", x"1FCF", x"1FD0", x"1FD1",
	x"1FD4", x"1FD5", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"1FD6", x"1FD7", x"1FD8", x"1FD9", x"1FDA", x"1FDB",
	x"1FDC", x"1FDD", x"1FDE", x"1FDF", x"1FE3", x"1FE4", x"1FE5", x"1FE6",
	x"1FE7", x"1FE8", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008",
	x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000"
	);

	-- Ask Xilinx synthesis to use block RAMs if possible
	attribute ram_style : string;
	attribute ram_style of RAM : signal is "block";
	-- Ask Quartus synthesis to use block RAMs if possible
	attribute ramstyle : string;
	attribute ramstyle of RAM : signal is "M10K";

begin
	p_RAM : process
	begin
		wait until rising_edge(I_MCKR);
		if I_En ='0' then
			if I_Wn = '0' then
				RAM(to_integer(unsigned(I_ADDR))) <= I_DATA;
			else
				O_DATA <= RAM(to_integer(unsigned(I_ADDR)));
			end if;
		end if;
	end process;
end RTL;