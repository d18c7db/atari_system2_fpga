--	(c) 2020 d18c7db(a)hotmail
--
--	This program is free software; you can redistribute it and/or modify it under
--	the terms of the GNU General Public License version 3 or, at your option,
--	any later version as published by the Free Software Foundation.
--
--	This program is distributed in the hope that it will be useful,
--	but WITHOUT ANY WARRANTY; without even the implied warranty of
--	MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.
--
-- For full details, see the GNU General Public License at www.gnu.org/licenses
--
-- generic 2K x 8 RAM definition

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;

entity RAM_2K8_0 is
	port(
		I_MCKR : in  std_logic;
		I_En   : in  std_logic;
		I_Wn   : in  std_logic;
		I_ADDR : in  std_logic_vector(10 downto 0);
		I_DATA : in  std_logic_vector( 7 downto 0);
		O_DATA : out std_logic_vector( 7 downto 0)
	);
end RAM_2K8_0;

architecture RTL of RAM_2K8_0 is
	type RAM_ARRAY_2Kx8 is array (0 to 2047) of std_logic_vector(7 downto 0);
	signal RAM : RAM_ARRAY_2Kx8 := (
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7",
	x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E1", x"EC", x"E7", x"E9", x"E9",
	x"EB", x"E8", x"00", x"DF", x"ED", x"DE", x"E6", x"E7", x"E1", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"00",
	x"00", x"00", x"39", x"71", x"64", x"2E", x"2A", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"3A", x"73", x"44", x"5E", x"2C", x"00", x"00", x"00", x"B0", x"AE", x"00", x"00", x"BA", x"00",
	x"BB", x"C1", x"00", x"C2", x"C4", x"00", x"00", x"00", x"00", x"00", x"00", x"E8", x"E7", x"E7", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B4", x"AF", x"B3", x"00", x"BD", x"B7",
	x"BC", x"C2", x"C7", x"C5", x"C7", x"CC", x"D0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"39", x"71", x"64", x"2E", x"2A", x"00", x"00", x"00", x"B7", x"B0", x"B4", x"00", x"C0", x"B8",
	x"BD", x"C3", x"C8", x"C8", x"CA", x"CD", x"D1", x"00", x"00", x"00", x"00", x"DF", x"E7", x"E5", x"00", x"00",
	x"00", x"00", x"3A", x"73", x"44", x"5E", x"2C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"C9", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"D9", x"D4", x"DA", x"DA", x"E2", x"E0", x"E6", x"EC", x"00", x"E7",
	x"FF", x"00", x"E5", x"00", x"E2", x"E1", x"EC", x"EB", x"EC", x"EB", x"DE", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"00",
	x"00", x"00", x"00", x"2A", x"4F", x"2A", x"79", x"42", x"53", x"32", x"00", x"59", x"2A", x"59", x"39", x"2E",
	x"2E", x"56", x"75", x"00", x"36", x"39", x"00", x"42", x"69", x"39", x"2E", x"60", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"2C", x"51", x"2C", x"7B", x"44", x"55", x"3D", x"00", x"5B", x"2C", x"5B", x"3A", x"5E",
	x"30", x"57", x"77", x"00", x"38", x"3A", x"4D", x"44", x"6B", x"3A", x"5E", x"62", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"DE", x"DF", x"DC", x"00", x"DE", x"EF", x"DC", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"E6", x"EC", x"DE", x"E2", x"EE", x"00", x"DA", x"DD", x"E5", x"EC", x"00", x"00", x"00", x"00",
	x"00", x"00", x"DA", x"E7", x"00", x"E8", x"E8", x"EC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"DB", x"DF", x"E5", x"EC", x"E9", x"E5", x"DC", x"7E", x"EB", x"EC", x"DD", x"E7", x"EC", x"00",
	x"00", x"00", x"E2", x"00", x"EE", x"E4", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"AD", x"AD", x"00", x"AD", x"00", x"00", x"A3", x"A3", x"A3", x"A3", x"A3", x"00", x"00",
	x"00", x"00", x"A3", x"A3", x"A3", x"A3", x"A3", x"A3", x"A3", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"A6", x"A4", x"A4", x"A6", x"A4", x"A6", x"00", x"A7", x"A5", x"A5", x"A7", x"A5", x"00", x"00",
	x"00", x"00", x"A7", x"A5", x"A5", x"A7", x"A5", x"A7", x"A5", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"A8", x"AA", x"A8", x"AA", x"A8", x"A8", x"00", x"AC", x"A9", x"A9", x"AC", x"A9", x"00", x"00",
	x"00", x"00", x"AC", x"A9", x"A9", x"AC", x"A9", x"AC", x"A9", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"A0", x"A0", x"A0", x"A2", x"A0", x"A2", x"00", x"A1", x"A1", x"A1", x"A3", x"A3", x"00", x"00",
	x"00", x"00", x"A1", x"A1", x"A1", x"A3", x"A3", x"A1", x"A1", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"A4", x"A4", x"A4", x"A6", x"A4", x"A6", x"00", x"A7", x"A5", x"A5", x"A7", x"A5", x"00", x"00",
	x"00", x"00", x"A7", x"A5", x"A5", x"A7", x"A5", x"A7", x"A5", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"A8", x"AA", x"A8", x"AA", x"A8", x"A8", x"00", x"AC", x"A9", x"A9", x"AC", x"A9", x"00", x"00",
	x"00", x"00", x"AC", x"A9", x"A9", x"AC", x"A9", x"AC", x"A9", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"A2", x"A0", x"A0", x"A2", x"A0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"A1", x"A1", x"A1", x"A3", x"A3", x"A3", x"A3", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"A6", x"A4", x"A4", x"A6", x"A4", x"00", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"00",
	x"00", x"00", x"A7", x"A5", x"A5", x"A7", x"A5", x"A7", x"A5", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"A8", x"AA", x"A8", x"AA", x"A8", x"00", x"E1", x"EB", x"00", x"DA", x"DE", x"DB", x"F2", x"00",
	x"00", x"00", x"AC", x"A9", x"A9", x"AC", x"A9", x"AC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"A2", x"A0", x"A0", x"A2", x"A0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"A6", x"A4", x"A4", x"A6", x"A4", x"00", x"EC", x"E8", x"EC", x"ED", x"E2", x"DF", x"00", x"00",
	x"00", x"00", x"00", x"FA", x"FA", x"FA", x"FA", x"FA", x"00", x"F9", x"A1", x"A1", x"A1", x"A3", x"A1", x"A1",
	x"A1", x"F9", x"A8", x"AA", x"A8", x"AA", x"A8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"F9", x"A7", x"A7", x"A7", x"A7", x"A7", x"A7",
	x"A7", x"F9", x"A0", x"A0", x"A0", x"A2", x"A0", x"00", x"00", x"AD", x"AD", x"00", x"AD", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FB", x"A4", x"A4", x"A4", x"A6", x"A4", x"00", x"A6", x"A4", x"A4", x"A6", x"A4", x"A6", x"00", x"00",
	x"00", x"00", x"DA", x"E7", x"EB", x"E7", x"DE", x"85", x"E9", x"F8", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"A8", x"AA", x"A8", x"AA", x"A8", x"00", x"A8", x"AA", x"A8", x"AA", x"A8", x"A8", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F9", x"E2", x"A1", x"00", x"00", x"E8", x"E0",
	x"00", x"00", x"A2", x"A0", x"A0", x"A2", x"A0", x"00", x"A0", x"A0", x"A0", x"A2", x"A0", x"A2", x"00", x"00",
	x"00", x"00", x"F0", x"EB", x"EC", x"00", x"00", x"00", x"00", x"F9", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"A6", x"A4", x"A4", x"A6", x"A4", x"00", x"A4", x"A4", x"A4", x"A6", x"A4", x"A6", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F9", x"E8", x"7E", x"DB", x"ED", x"FF", x"A2",
	x"00", x"00", x"A8", x"AA", x"A8", x"AA", x"A8", x"00", x"A8", x"AA", x"A8", x"AA", x"A8", x"A8", x"00", x"00",
	x"00", x"00", x"A3", x"A3", x"A3", x"A3", x"A3", x"A3", x"A3", x"F9", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"A0", x"A0", x"A0", x"A2", x"A0", x"00", x"A2", x"A0", x"A0", x"A2", x"A0", x"00", x"00", x"00",
	x"00", x"00", x"A7", x"A5", x"A5", x"A7", x"A5", x"A7", x"A5", x"F9", x"A3", x"A3", x"A3", x"A3", x"A3", x"A3",
	x"A3", x"00", x"A4", x"A4", x"A4", x"A6", x"A4", x"00", x"A6", x"A4", x"A4", x"A6", x"A4", x"A6", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
	);

	-- Ask Xilinx synthesis to use block RAMs if possible
	attribute ram_style : string;
	attribute ram_style of RAM : signal is "block";
	-- Ask Quartus synthesis to use block RAMs if possible
	attribute ramstyle : string;
	attribute ramstyle of RAM : signal is "M10K";

begin
	p_RAM : process
	begin
		wait until rising_edge(I_MCKR);
		if I_En ='0' then
			if I_Wn = '0' then
				RAM(to_integer(unsigned(I_ADDR))) <= I_DATA;
			else
				O_DATA <= RAM(to_integer(unsigned(I_ADDR)));
			end if;
		end if;
	end process;
end RTL;